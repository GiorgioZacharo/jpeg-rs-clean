`timescale 1 ns / 1 ps

module AESL_deadlock_detector (
    input reset,
    input clock);

    wire [1:0] proc_dep_vld_vec_0;
    reg [1:0] proc_dep_vld_vec_0_reg;
    wire [1:0] in_chan_dep_vld_vec_0;
    wire [5:0] in_chan_dep_data_vec_0;
    wire [1:0] token_in_vec_0;
    wire [1:0] out_chan_dep_vld_vec_0;
    wire [2:0] out_chan_dep_data_0;
    wire [1:0] token_out_vec_0;
    wire dl_detect_out_0;
    wire dep_chan_vld_1_0;
    wire [2:0] dep_chan_data_1_0;
    wire token_1_0;
    wire dep_chan_vld_2_0;
    wire [2:0] dep_chan_data_2_0;
    wire token_2_0;
    wire [1:0] proc_dep_vld_vec_1;
    reg [1:0] proc_dep_vld_vec_1_reg;
    wire [1:0] in_chan_dep_vld_vec_1;
    wire [5:0] in_chan_dep_data_vec_1;
    wire [1:0] token_in_vec_1;
    wire [1:0] out_chan_dep_vld_vec_1;
    wire [2:0] out_chan_dep_data_1;
    wire [1:0] token_out_vec_1;
    wire dl_detect_out_1;
    wire dep_chan_vld_0_1;
    wire [2:0] dep_chan_data_0_1;
    wire token_0_1;
    wire dep_chan_vld_2_1;
    wire [2:0] dep_chan_data_2_1;
    wire token_2_1;
    wire [1:0] proc_dep_vld_vec_2;
    reg [1:0] proc_dep_vld_vec_2_reg;
    wire [1:0] in_chan_dep_vld_vec_2;
    wire [5:0] in_chan_dep_data_vec_2;
    wire [1:0] token_in_vec_2;
    wire [1:0] out_chan_dep_vld_vec_2;
    wire [2:0] out_chan_dep_data_2;
    wire [1:0] token_out_vec_2;
    wire dl_detect_out_2;
    wire dep_chan_vld_0_2;
    wire [2:0] dep_chan_data_0_2;
    wire token_0_2;
    wire dep_chan_vld_1_2;
    wire [2:0] dep_chan_data_1_2;
    wire token_1_2;
    wire [2:0] dl_in_vec;
    wire dl_detect_out;
    wire [2:0] origin;
    wire token_clear;

    reg ap_done_reg_0;
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            ap_done_reg_0 <= 'b0;
        end
        else begin
            ap_done_reg_0 <= AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.Loop_0_proc19_U0.ap_done;
        end
    end

    reg ap_done_reg_1;
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            ap_done_reg_1 <= 'b0;
        end
        else begin
            ap_done_reg_1 <= AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.Loop_1_proc_U0.ap_done;
        end
    end

    reg ap_done_reg_2;
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            ap_done_reg_2 <= 'b0;
        end
        else begin
            ap_done_reg_2 <= AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.memcpy_omatrix_out_b_U0.ap_done;
        end
    end

    // delay ap_idle for one cycle
    reg [0:0] AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd$dataflow_in_loop_U0$Loop_0_proc19_U0$ap_idle;
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd$dataflow_in_loop_U0$Loop_0_proc19_U0$ap_idle <= 'b0;
        end
        else begin
            AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd$dataflow_in_loop_U0$Loop_0_proc19_U0$ap_idle <= AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.Loop_0_proc19_U0.ap_idle;
        end
    end
    // Process: AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.Loop_0_proc19_U0
    AESL_deadlock_detect_unit #(3, 0, 2, 2) AESL_deadlock_detect_unit_0 (
        .reset(reset),
        .clock(clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_0),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_0),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_0),
        .token_in_vec(token_in_vec_0),
        .dl_detect_in(dl_detect_out),
        .origin(origin[0]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_0),
        .out_chan_dep_data(out_chan_dep_data_0),
        .token_out_vec(token_out_vec_0),
        .dl_detect_out(dl_in_vec[0]));

    assign proc_dep_vld_vec_0[0] = dl_detect_out ? proc_dep_vld_vec_0_reg[0] : (~AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.in1_buf_0_U.i_full_n & AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.Loop_0_proc19_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.in1_buf_0_U.t_read | ~AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.in1_buf_1_U.i_full_n & AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.Loop_0_proc19_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.in1_buf_1_U.t_read | ~AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.in1_buf_2_U.i_full_n & AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.Loop_0_proc19_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.in1_buf_2_U.t_read | ~AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.in1_buf_3_U.i_full_n & AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.Loop_0_proc19_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.in1_buf_3_U.t_read | ~AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.in1_buf_4_U.i_full_n & AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.Loop_0_proc19_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.in1_buf_4_U.t_read | ~AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.in1_buf_5_U.i_full_n & AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.Loop_0_proc19_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.in1_buf_5_U.t_read | ~AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.in1_buf_6_U.i_full_n & AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.Loop_0_proc19_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.in1_buf_6_U.t_read | ~AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.in1_buf_7_U.i_full_n & AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.Loop_0_proc19_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.in1_buf_7_U.t_read | ~AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.in1_buf_8_U.i_full_n & AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.Loop_0_proc19_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.in1_buf_8_U.t_read | ~AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.in1_buf_9_U.i_full_n & AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.Loop_0_proc19_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.in1_buf_9_U.t_read | ~AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.in1_buf_10_U.i_full_n & AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.Loop_0_proc19_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.in1_buf_10_U.t_read | ~AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.in1_buf_11_U.i_full_n & AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.Loop_0_proc19_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.in1_buf_11_U.t_read | ~AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.in1_buf_12_U.i_full_n & AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.Loop_0_proc19_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.in1_buf_12_U.t_read | ~AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.in1_buf_13_U.i_full_n & AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.Loop_0_proc19_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.in1_buf_13_U.t_read | ~AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.in1_buf_14_U.i_full_n & AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.Loop_0_proc19_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.in1_buf_14_U.t_read | ~AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.in1_buf_15_U.i_full_n & AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.Loop_0_proc19_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.in1_buf_15_U.t_read | ~AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.Loop_0_proc19_U0.imatrix_offset_out_blk_n);
    assign proc_dep_vld_vec_0[1] = dl_detect_out ? proc_dep_vld_vec_0_reg[1] : (~AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.Loop_0_proc19_U0.i_0_i_i_c_blk_n | ~AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.Loop_0_proc19_U0.omatrix_offset_out_blk_n);
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            proc_dep_vld_vec_0_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_0_reg <= proc_dep_vld_vec_0;
        end
    end
    assign in_chan_dep_vld_vec_0[0] = dep_chan_vld_1_0;
    assign in_chan_dep_data_vec_0[2 : 0] = dep_chan_data_1_0;
    assign token_in_vec_0[0] = token_1_0;
    assign in_chan_dep_vld_vec_0[1] = dep_chan_vld_2_0;
    assign in_chan_dep_data_vec_0[5 : 3] = dep_chan_data_2_0;
    assign token_in_vec_0[1] = token_2_0;
    assign dep_chan_vld_0_1 = out_chan_dep_vld_vec_0[0];
    assign dep_chan_data_0_1 = out_chan_dep_data_0;
    assign token_0_1 = token_out_vec_0[0];
    assign dep_chan_vld_0_2 = out_chan_dep_vld_vec_0[1];
    assign dep_chan_data_0_2 = out_chan_dep_data_0;
    assign token_0_2 = token_out_vec_0[1];

    // delay ap_idle for one cycle
    reg [0:0] AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd$dataflow_in_loop_U0$Loop_1_proc_U0$ap_idle;
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd$dataflow_in_loop_U0$Loop_1_proc_U0$ap_idle <= 'b0;
        end
        else begin
            AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd$dataflow_in_loop_U0$Loop_1_proc_U0$ap_idle <= AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.Loop_1_proc_U0.ap_idle;
        end
    end
    // Process: AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.Loop_1_proc_U0
    AESL_deadlock_detect_unit #(3, 1, 2, 2) AESL_deadlock_detect_unit_1 (
        .reset(reset),
        .clock(clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_1),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_1),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_1),
        .token_in_vec(token_in_vec_1),
        .dl_detect_in(dl_detect_out),
        .origin(origin[1]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_1),
        .out_chan_dep_data(out_chan_dep_data_1),
        .token_out_vec(token_out_vec_1),
        .dl_detect_out(dl_in_vec[1]));

    assign proc_dep_vld_vec_1[0] = dl_detect_out ? proc_dep_vld_vec_1_reg[0] : (~AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.in1_buf_0_U.t_empty_n & (AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.Loop_1_proc_U0.ap_ready | AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.Loop_1_proc_U0.ap_idle) & ~AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.in1_buf_0_U.i_write | ~AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.Loop_1_proc_U0.imatrix_offset_blk_n | ~AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.in1_buf_1_U.t_empty_n & (AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.Loop_1_proc_U0.ap_ready | AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.Loop_1_proc_U0.ap_idle) & ~AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.in1_buf_1_U.i_write | ~AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.in1_buf_2_U.t_empty_n & (AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.Loop_1_proc_U0.ap_ready | AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.Loop_1_proc_U0.ap_idle) & ~AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.in1_buf_2_U.i_write | ~AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.in1_buf_3_U.t_empty_n & (AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.Loop_1_proc_U0.ap_ready | AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.Loop_1_proc_U0.ap_idle) & ~AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.in1_buf_3_U.i_write | ~AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.in1_buf_4_U.t_empty_n & (AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.Loop_1_proc_U0.ap_ready | AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.Loop_1_proc_U0.ap_idle) & ~AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.in1_buf_4_U.i_write | ~AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.in1_buf_5_U.t_empty_n & (AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.Loop_1_proc_U0.ap_ready | AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.Loop_1_proc_U0.ap_idle) & ~AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.in1_buf_5_U.i_write | ~AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.in1_buf_6_U.t_empty_n & (AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.Loop_1_proc_U0.ap_ready | AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.Loop_1_proc_U0.ap_idle) & ~AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.in1_buf_6_U.i_write | ~AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.in1_buf_7_U.t_empty_n & (AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.Loop_1_proc_U0.ap_ready | AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.Loop_1_proc_U0.ap_idle) & ~AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.in1_buf_7_U.i_write | ~AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.in1_buf_8_U.t_empty_n & (AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.Loop_1_proc_U0.ap_ready | AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.Loop_1_proc_U0.ap_idle) & ~AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.in1_buf_8_U.i_write | ~AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.in1_buf_9_U.t_empty_n & (AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.Loop_1_proc_U0.ap_ready | AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.Loop_1_proc_U0.ap_idle) & ~AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.in1_buf_9_U.i_write | ~AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.in1_buf_10_U.t_empty_n & (AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.Loop_1_proc_U0.ap_ready | AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.Loop_1_proc_U0.ap_idle) & ~AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.in1_buf_10_U.i_write | ~AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.in1_buf_11_U.t_empty_n & (AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.Loop_1_proc_U0.ap_ready | AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.Loop_1_proc_U0.ap_idle) & ~AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.in1_buf_11_U.i_write | ~AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.in1_buf_12_U.t_empty_n & (AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.Loop_1_proc_U0.ap_ready | AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.Loop_1_proc_U0.ap_idle) & ~AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.in1_buf_12_U.i_write | ~AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.in1_buf_13_U.t_empty_n & (AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.Loop_1_proc_U0.ap_ready | AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.Loop_1_proc_U0.ap_idle) & ~AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.in1_buf_13_U.i_write | ~AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.in1_buf_14_U.t_empty_n & (AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.Loop_1_proc_U0.ap_ready | AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.Loop_1_proc_U0.ap_idle) & ~AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.in1_buf_14_U.i_write | ~AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.in1_buf_15_U.t_empty_n & (AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.Loop_1_proc_U0.ap_ready | AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.Loop_1_proc_U0.ap_idle) & ~AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.in1_buf_15_U.i_write);
    assign proc_dep_vld_vec_1[1] = dl_detect_out ? proc_dep_vld_vec_1_reg[1] : (~AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.out_buf_0_U.i_full_n & AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.Loop_1_proc_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.out_buf_0_U.t_read | ~AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.out_buf_1_U.i_full_n & AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.Loop_1_proc_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.out_buf_1_U.t_read | ~AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.out_buf_2_U.i_full_n & AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.Loop_1_proc_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.out_buf_2_U.t_read | ~AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.out_buf_3_U.i_full_n & AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.Loop_1_proc_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.out_buf_3_U.t_read | ~AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.out_buf_4_U.i_full_n & AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.Loop_1_proc_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.out_buf_4_U.t_read | ~AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.out_buf_5_U.i_full_n & AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.Loop_1_proc_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.out_buf_5_U.t_read | ~AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.out_buf_6_U.i_full_n & AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.Loop_1_proc_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.out_buf_6_U.t_read | ~AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.out_buf_7_U.i_full_n & AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.Loop_1_proc_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.out_buf_7_U.t_read | ~AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.out_buf_8_U.i_full_n & AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.Loop_1_proc_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.out_buf_8_U.t_read | ~AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.out_buf_9_U.i_full_n & AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.Loop_1_proc_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.out_buf_9_U.t_read | ~AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.out_buf_10_U.i_full_n & AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.Loop_1_proc_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.out_buf_10_U.t_read | ~AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.out_buf_11_U.i_full_n & AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.Loop_1_proc_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.out_buf_11_U.t_read | ~AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.out_buf_12_U.i_full_n & AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.Loop_1_proc_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.out_buf_12_U.t_read | ~AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.out_buf_13_U.i_full_n & AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.Loop_1_proc_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.out_buf_13_U.t_read | ~AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.out_buf_14_U.i_full_n & AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.Loop_1_proc_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.out_buf_14_U.t_read | ~AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.out_buf_15_U.i_full_n & AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.Loop_1_proc_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.out_buf_15_U.t_read);
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            proc_dep_vld_vec_1_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_1_reg <= proc_dep_vld_vec_1;
        end
    end
    assign in_chan_dep_vld_vec_1[0] = dep_chan_vld_0_1;
    assign in_chan_dep_data_vec_1[2 : 0] = dep_chan_data_0_1;
    assign token_in_vec_1[0] = token_0_1;
    assign in_chan_dep_vld_vec_1[1] = dep_chan_vld_2_1;
    assign in_chan_dep_data_vec_1[5 : 3] = dep_chan_data_2_1;
    assign token_in_vec_1[1] = token_2_1;
    assign dep_chan_vld_1_0 = out_chan_dep_vld_vec_1[0];
    assign dep_chan_data_1_0 = out_chan_dep_data_1;
    assign token_1_0 = token_out_vec_1[0];
    assign dep_chan_vld_1_2 = out_chan_dep_vld_vec_1[1];
    assign dep_chan_data_1_2 = out_chan_dep_data_1;
    assign token_1_2 = token_out_vec_1[1];

    // delay ap_idle for one cycle
    reg [0:0] AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd$dataflow_in_loop_U0$memcpy_omatrix_out_b_U0$ap_idle;
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd$dataflow_in_loop_U0$memcpy_omatrix_out_b_U0$ap_idle <= 'b0;
        end
        else begin
            AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd$dataflow_in_loop_U0$memcpy_omatrix_out_b_U0$ap_idle <= AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.memcpy_omatrix_out_b_U0.ap_idle;
        end
    end
    // Process: AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.memcpy_omatrix_out_b_U0
    AESL_deadlock_detect_unit #(3, 2, 2, 2) AESL_deadlock_detect_unit_2 (
        .reset(reset),
        .clock(clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_2),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_2),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_2),
        .token_in_vec(token_in_vec_2),
        .dl_detect_in(dl_detect_out),
        .origin(origin[2]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_2),
        .out_chan_dep_data(out_chan_dep_data_2),
        .token_out_vec(token_out_vec_2),
        .dl_detect_out(dl_in_vec[2]));

    assign proc_dep_vld_vec_2[0] = dl_detect_out ? proc_dep_vld_vec_2_reg[0] : (~AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.memcpy_omatrix_out_b_U0.omatrix_offset_blk_n | ~AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.memcpy_omatrix_out_b_U0.i_0_i_i_c_blk_n);
    assign proc_dep_vld_vec_2[1] = dl_detect_out ? proc_dep_vld_vec_2_reg[1] : (~AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.out_buf_0_U.t_empty_n & (AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.memcpy_omatrix_out_b_U0.ap_ready | AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.memcpy_omatrix_out_b_U0.ap_idle) & ~AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.out_buf_0_U.i_write | ~AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.out_buf_1_U.t_empty_n & (AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.memcpy_omatrix_out_b_U0.ap_ready | AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.memcpy_omatrix_out_b_U0.ap_idle) & ~AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.out_buf_1_U.i_write | ~AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.out_buf_2_U.t_empty_n & (AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.memcpy_omatrix_out_b_U0.ap_ready | AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.memcpy_omatrix_out_b_U0.ap_idle) & ~AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.out_buf_2_U.i_write | ~AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.out_buf_3_U.t_empty_n & (AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.memcpy_omatrix_out_b_U0.ap_ready | AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.memcpy_omatrix_out_b_U0.ap_idle) & ~AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.out_buf_3_U.i_write | ~AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.out_buf_4_U.t_empty_n & (AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.memcpy_omatrix_out_b_U0.ap_ready | AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.memcpy_omatrix_out_b_U0.ap_idle) & ~AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.out_buf_4_U.i_write | ~AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.out_buf_5_U.t_empty_n & (AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.memcpy_omatrix_out_b_U0.ap_ready | AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.memcpy_omatrix_out_b_U0.ap_idle) & ~AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.out_buf_5_U.i_write | ~AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.out_buf_6_U.t_empty_n & (AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.memcpy_omatrix_out_b_U0.ap_ready | AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.memcpy_omatrix_out_b_U0.ap_idle) & ~AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.out_buf_6_U.i_write | ~AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.out_buf_7_U.t_empty_n & (AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.memcpy_omatrix_out_b_U0.ap_ready | AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.memcpy_omatrix_out_b_U0.ap_idle) & ~AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.out_buf_7_U.i_write | ~AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.out_buf_8_U.t_empty_n & (AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.memcpy_omatrix_out_b_U0.ap_ready | AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.memcpy_omatrix_out_b_U0.ap_idle) & ~AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.out_buf_8_U.i_write | ~AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.out_buf_9_U.t_empty_n & (AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.memcpy_omatrix_out_b_U0.ap_ready | AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.memcpy_omatrix_out_b_U0.ap_idle) & ~AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.out_buf_9_U.i_write | ~AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.out_buf_10_U.t_empty_n & (AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.memcpy_omatrix_out_b_U0.ap_ready | AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.memcpy_omatrix_out_b_U0.ap_idle) & ~AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.out_buf_10_U.i_write | ~AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.out_buf_11_U.t_empty_n & (AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.memcpy_omatrix_out_b_U0.ap_ready | AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.memcpy_omatrix_out_b_U0.ap_idle) & ~AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.out_buf_11_U.i_write | ~AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.out_buf_12_U.t_empty_n & (AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.memcpy_omatrix_out_b_U0.ap_ready | AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.memcpy_omatrix_out_b_U0.ap_idle) & ~AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.out_buf_12_U.i_write | ~AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.out_buf_13_U.t_empty_n & (AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.memcpy_omatrix_out_b_U0.ap_ready | AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.memcpy_omatrix_out_b_U0.ap_idle) & ~AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.out_buf_13_U.i_write | ~AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.out_buf_14_U.t_empty_n & (AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.memcpy_omatrix_out_b_U0.ap_ready | AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.memcpy_omatrix_out_b_U0.ap_idle) & ~AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.out_buf_14_U.i_write | ~AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.out_buf_15_U.t_empty_n & (AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.memcpy_omatrix_out_b_U0.ap_ready | AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.memcpy_omatrix_out_b_U0.ap_idle) & ~AESL_inst_IZigzagMatrix_f2r_forBody_s2e_forEnd.dataflow_in_loop_U0.out_buf_15_U.i_write);
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            proc_dep_vld_vec_2_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_2_reg <= proc_dep_vld_vec_2;
        end
    end
    assign in_chan_dep_vld_vec_2[0] = dep_chan_vld_0_2;
    assign in_chan_dep_data_vec_2[2 : 0] = dep_chan_data_0_2;
    assign token_in_vec_2[0] = token_0_2;
    assign in_chan_dep_vld_vec_2[1] = dep_chan_vld_1_2;
    assign in_chan_dep_data_vec_2[5 : 3] = dep_chan_data_1_2;
    assign token_in_vec_2[1] = token_1_2;
    assign dep_chan_vld_2_0 = out_chan_dep_vld_vec_2[0];
    assign dep_chan_data_2_0 = out_chan_dep_data_2;
    assign token_2_0 = token_out_vec_2[0];
    assign dep_chan_vld_2_1 = out_chan_dep_vld_vec_2[1];
    assign dep_chan_data_2_1 = out_chan_dep_data_2;
    assign token_2_1 = token_out_vec_2[1];


    AESL_deadlock_report_unit #(3) AESL_deadlock_report_unit_inst (
        .reset(reset),
        .clock(clock),
        .dl_in_vec(dl_in_vec),
        .dl_detect_out(dl_detect_out),
        .origin(origin),
        .token_clear(token_clear));

endmodule
